library verilog;
use verilog.vl_types.all;
entity BLOCO_PRINCIPAL_vlg_vec_tst is
end BLOCO_PRINCIPAL_vlg_vec_tst;
