LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- ESTA SEGUNDA IMPLEMENTAÇÃO SERA COM BASE NO FSM PARA VHDL, DEMONSTRAD POR VOLNEI

ENTITY COUNTER_MOD5_V2 IS
	PORT(
			R : IN STD_LOGIC;
			CLK : IN STD_LOGIC;
			QOUT : OUT STD_LOGIC_VECTOR( 2 DOWNTO 0)
			);
	
END COUNTER_MOD5_V2;

ARCHITECTURE LOGIC OF COUNTER_MOD5_V2 IS

TYPE LIST_STATES IS (ZERO, UM, DOIS, TRES, QUATRO);
SIGNAL PR_STATE, NX_STATE : LIST_STATES;

BEGIN

-- BLOCO COMBINACIONAL: PROCESSANDO
-- PR_STATE E PRODUZINDO NX_STATE E A SAIDA

-- SEMPRE QUE PR_STATE SOFRE ALTERAÇÕES, ESTE BLOCO
-- ENTRA EM EXECUÇÃO
PROCESS( PR_STATE )
BEGIN



	-- PARA CADA ESTADO, DEFINA A SAIDA E O NX_STATE
	CASE PR_STATE IS
	
		WHEN ZERO =>
		
			QOUT <= "000";

			NX_STATE <= UM;
			
		WHEN UM =>
		
			QOUT <= "001";

			NX_STATE <= DOIS;
			
		WHEN DOIS =>
			
			QOUT <= "010";

			NX_STATE <= TRES;
			
		WHEN TRES =>
		
			QOUT <= "011";

			NX_STATE <= QUATRO;
			
		WHEN QUATRO =>
		
			QOUT <= "100";

			NX_STATE <= ZERO;
			
	END CASE;
END PROCESS;
	
-- BLOCO SEQUENCIAL: CARREGA O NX_STATE PARA
-- PR_STATE

	PROCESS( CLK , R )
	BEGIN
	
		IF( R = '1') THEN
			PR_STATE <= ZERO;
		ELSIF( FALLING_EDGE(CLK) ) THEN
			PR_STATE <= NX_STATE;
		END IF;
	END PROCESS;

END LOGIC;