LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;

ENTITY SELETOR_FREQUENCIA IS
PORT(
		CLK_IN : IN STD_LOGIC;
		CLK_ALT : IN STD_LOGIC;
		COMANDO : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		CLK_OUT : OUT STD_LOGIC
	);
END SELETOR_FREQUENCIA;

ARCHITECTURE LOGICA OF SELETOR_FREQUENCIA IS

SIGNAL CONSTANTE : STD_LOGIC := '1';
SIGNAL CLOCK_1HZ : STD_LOGIC := '1';
SIGNAL CLOCK_nHZ : STD_LOGIC := '1';

BEGIN

PROCESS(CLK_IN)
	VARIABLE COUNT : INTEGER := 1;
	VARIABLE N : INTEGER := 1;
BEGIN
	IF( CLK_IN'EVENT AND CLK_IN = '0') THEN
		COUNT:= COUNT +1;
		
		IF(COUNT = 13500000) THEN
			CLOCK_1HZ <= NOT CLOCK_1HZ;
			
			
		END IF;
		-- 2Hz = 675000
		-- 4Hz = 337500
		-- 8Hz = 168750
		IF(COUNT = N*675000) THEN
			
			CLOCK_nHZ <= NOT CLOCK_nHZ;
			N := N + 1;
			
			IF(COUNT = 13500000) THEN
				N := 1;
				COUNT := 1;
			END IF;
		END IF;
	END IF;
END PROCESS;

-- MULTIPLEXAÇÃO DO CLOCK

WITH COMANDO SELECT
CLK_OUT <=   CLK_ALT WHEN "00",
			  CLOCK_1HZ WHEN "01",
			  CLOCK_nHZ WHEN "10",
			  CONSTANTE WHEN "11";
				
END LOGICA;