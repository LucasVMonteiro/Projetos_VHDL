library verilog;
use verilog.vl_types.all;
entity CONVERSOR_1KHZ_vlg_sample_tst is
    port(
        CLK_I           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end CONVERSOR_1KHZ_vlg_sample_tst;
