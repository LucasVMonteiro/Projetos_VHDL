LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
-- CODIGO PREPARADO PARA CLOCK DE 50MHz

ENTITY BLOCO_PRINCIPAL IS
PORT(

		CLK_IN : IN STD_LOGIC;
		MONITOR_CLOCK_RED : OUT STD_LOGIC;
		MONITOR_CLOCK_1S : OUT STD_LOGIC;
		MONITOR_FLAG : OUT STD_LOGIC;
		MONITOR_ESPERA : OUT STD_LOGIC;
		SAIDA_RED : OUT STD_LOGIC_VECTOR( 17 DOWNTO 0)
		
		);
		
END BLOCO_PRINCIPAL;


ARCHITECTURE LOGICA OF BLOCO_PRINCIPAL IS

SIGNAL SINAL_CLK : STD_LOGIC:= '0';
CONSTANT FREQUENCIA : INTEGER := 50000000;
CONSTANT TEMPO : INTEGER := 10; -- EM SEGUNDOS
CONSTANT BITS_RED : INTEGER := 18;
--CONSTANT BITS_GREEN : INTEGER := 8;
CONSTANT MEIO_PERIODO_BIT_RED : INTEGER := 1000000*TEMPO/(2*BITS_RED);
CONSTANT PULSOS_MEIO_PERIODO_BIT_RED : INTEGER := MEIO_PERIODO_BIT_RED*(FREQUENCIA/1000000);
SIGNAL CLOCK_RED : STD_LOGIC := '0';

SIGNAL LEDS_R : STD_LOGIC_VECTOR(17 DOWNTO 0):= "111111111111111111";
SIGNAL CLOCK_1S : STD_LOGIC := '0';
SIGNAL BITS_R_DESLOCADOS_PROCESS_CLOCK_RED : INTEGER := 0;
SIGNAL ESPERA_R : STD_LOGIC := '0';

BEGIN

PROCESS(CLK_IN)
	VARIABLE CONTADOR_SEGUNDOS : INTEGER := 1;
	VARIABLE CONTADOR_CLOCK_RED : INTEGER := 1;
	VARIABLE BITS_R_DESLOCADOS : INTEGER := 0;
	

BEGIN


	IF( FALLING_EDGE(CLK_IN) ) THEN
		CONTADOR_SEGUNDOS := CONTADOR_SEGUNDOS + 1;
		IF( ESPERA_R = '0') THEN
			CONTADOR_CLOCK_RED := CONTADOR_CLOCK_RED + 1;	
		END IF;
		
		IF( CONTADOR_CLOCK_RED = PULSOS_MEIO_PERIODO_BIT_RED AND ESPERA_R = '0') THEN
			-- O TOTAL DE BITS RED DESLOCADOS ATINGIU O VALOR MAXIMO E O CONTADOR DE SEGUNDOS NÃO? ENTAO FAÇA
			IF ( BITS_R_DESLOCADOS = BITS_RED AND CLOCK_RED = '1' AND CONTADOR_SEGUNDOS < TEMPO*FREQUENCIA ) THEN
				BITS_R_DESLOCADOS := 0;
				ESPERA_R <= '1';
				-- SINALIZE PARA QUE INICIE O CONTADOR GREEN
				
			-- SE NAO, APENAS O TOTAL DE BITS RED DESLOCADOS ATINGIU O VALOR MAXIMO? ENTAO FAÇA
			ELSIF( BITS_R_DESLOCADOS = BITS_RED ) THEN
				BITS_R_DESLOCADOS := 0;
			
			-- SE NENHUM DOS CASOS ANTERIORES, ENTAO...
			ELSE
				BITS_R_DESLOCADOS := BITS_R_DESLOCADOS_PROCESS_CLOCK_RED;
				CLOCK_RED <= NOT CLOCK_RED;
				
			END IF;
			CONTADOR_CLOCK_RED := 1;
		END IF;
		-- CONTAR ATE "FREQUENCIA" LEVA 1 SEGUNDO
		-- CONTAR ATE "N*FREQUENCIA" LEVA N SEGUNDOS
		IF( CONTADOR_SEGUNDOS = TEMPO*FREQUENCIA ) THEN
			CONTADOR_SEGUNDOS := 0;
			ESPERA_R <= '0';
			CLOCK_1S <= NOT CLOCK_1S;
			
		END IF;
	END IF;
END PROCESS;
MONITOR_CLOCK_RED <= CLOCK_RED;
MONITOR_CLOCK_1S  <= CLOCK_1S;
MONITOR_ESPERA    <= ESPERA_R;
--MONITOR_FLAG      <= 
PROCESS(CLOCK_RED)
BEGIN
	IF( FALLING_EDGE(CLOCK_RED) )THEN 
		LEDS_R <= STD_LOGIC_VECTOR(SHIFT_RIGHT(UNSIGNED(LEDS_R),1));
		
		IF( BITS_R_DESLOCADOS_PROCESS_CLOCK_RED = BITS_RED) THEN
			BITS_R_DESLOCADOS_PROCESS_CLOCK_RED <= 0;
			
		ELSE 
			BITS_R_DESLOCADOS_PROCESS_CLOCK_RED <= BITS_R_DESLOCADOS_PROCESS_CLOCK_RED + 1;
		
		END IF;
		IF ( LEDS_R = "000000000000000000" AND ESPERA_R = '0') THEN
			LEDS_R <= "111111111111111111";
		END IF;
		
	END IF;
END PROCESS;

SAIDA_RED <= LEDS_R;
END LOGICA;