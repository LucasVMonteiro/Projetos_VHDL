library verilog;
use verilog.vl_types.all;
entity CONVERSOR_1KHZ is
    port(
        CLK_I           : in     vl_logic;
        CLK_O           : out    vl_logic
    );
end CONVERSOR_1KHZ;
