LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL; -- REFERENTE AO COMANDO UNSIGNED; VER CAPITULO 11 DE 'VHDL DECRICAO E SINTESE DE CIRCUITOS DIGITASI' d'AMORE

ENTITY BLOCO_CONTADOR23 IS
	PORT(
			CLK_IN : IN STD_LOGIC;
		
			-- UTILIZAR SAIDAS DE 7BITS PARA UM DECODIFICADOR DE 7 SEGMENTOS 
			-- 7 DOWNTO 0     ->   MSB / 7 / 6 / 5 / 4 / 3 / 2 / 1 / 0 / LSB
			-- 0 TO 7     ->    	  LSB / 0 / 1 / 2 / 3 / 4 / 5 / 6 / 7 / MSB
 			SAIDA : OUT STD_LOGIC_VECTOR( 7 DOWNTO 0)
	
	);
END BLOCO_CONTADOR23;

ARCHITECTURE LOGIC OF BLOCO_CONTADOR23 IS
BEGIN
-- PORQUE UTILIZAR UNSIGNED EM: ACUMULADOR_A := STD_LOGIC_VECTOR( UNSIGNED(ACUMULADOR_A) + "0001");?
-- RESPOSTA: OPERAÇÃO DE SOMA + COM VETORES PRECISA TER EXPLICITADO SE 
-- O VETOR BINARIO POSSUI BIT DE SINAL(SIGNED) OU NAO POSSUI( UNSIGNED)

PROCESSO_CONTADOR: PROCESS(CLK_IN)
		VARIABLE ACUMULADOR_UNIDADE: STD_LOGIC_VECTOR( 3 DOWNTO 0 );
		VARIABLE ACUMULADOR_DEZENA: STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	BEGIN

		IF ( CLK_IN'EVENT AND CLK_IN = '0' ) THEN 
		
			IF ( ACUMULADOR_UNIDADE >= "1001") THEN -- SE X9
				ACUMULADOR_UNIDADE := "0000";
				ACUMULADOR_DEZENA := STD_LOGIC_VECTOR( UNSIGNED(ACUMULADOR_DEZENA) + "0001");
				
			ELSIF( ACUMULADOR_DEZENA >= "0010" AND ACUMULADOR_UNIDADE >= "0011") THEN -- SE 23
			
				ACUMULADOR_UNIDADE := "0000";
				ACUMULADOR_DEZENA := "0000";

			ELSE
				ACUMULADOR_UNIDADE := STD_LOGIC_VECTOR( UNSIGNED(ACUMULADOR_UNIDADE) + "0001");
				
			END IF;
		END IF;
		
		
		
		SAIDA <=  ACUMULADOR_DEZENA & ACUMULADOR_UNIDADE;
	END PROCESS PROCESSO_CONTADOR;

END LOGIC;