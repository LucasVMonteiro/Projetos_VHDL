library verilog;
use verilog.vl_types.all;
entity FSM_MEALY_1_vlg_vec_tst is
end FSM_MEALY_1_vlg_vec_tst;
