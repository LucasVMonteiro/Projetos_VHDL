library verilog;
use verilog.vl_types.all;
entity COUNTER_MOD5_V1_vlg_vec_tst is
end COUNTER_MOD5_V1_vlg_vec_tst;
