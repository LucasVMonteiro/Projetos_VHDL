LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- ESTA PRIMEIR IMPLEMENTAÇÃO SERA COM BASE NO CIRCUITO LOGICO MONTADO

ENTITY COUNTER_MOD5_V1 IS
	PORT(
			R : IN STD_LOGIC;
			CLK : IN STD_LOGIC;
			QOUT : OUT STD_LOGIC_VECTOR( 2 DOWNTO 0)
			);
	
END COUNTER_MOD5_V1;

ARCHITECTURE LOGIC OF COUNTER_MOD5_V1 IS

SIGNAL D2, D1, D0 : STD_LOGIC := '0';
SIGNAL Q2, Q1, Q0 : STD_LOGIC := '0';

BEGIN
-- COMPORTAMENTO DOS 3 FF

PROCESS( CLK, R)
BEGIN
	IF FALLING_EDGE(CLK) THEN
		Q2 <= D2;
		Q1 <= D1;
		Q0 <= D0;
	END IF;
END PROCESS;

D0 <= (NOT Q0) AND (NOT Q2) AND (NOT R);
D1 <= ( Q1 AND (NOT Q0) AND (NOT R)) OR ( Q0 AND (NOT Q1) AND (NOT R));
D2 <= Q1 AND Q0 AND (NOT R);

QOUT <= Q2 & Q1 & Q0;

END LOGIC;