LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-- ESSE MODULO CONVERTE 27MHZ EM 1KHZ

-- PERIODO FUNDAMENTAL DE 1KHZ = 1/1000 = 0.001s

-- CLOCK FPGA 27MHZ = 27_000_000 CICLOS/S
-- ENTAO 	 1s => 27000000
-- 	   0.001s => 0.001  X 27000000 = 27000
--      0.0005s => 0.0005 X 27000000 = 13500
--
-- AO CONTAR 13500 CICLOS, PASSA-SE 0.0005s
-- E ALTERNANDO O SINAL DE CLK NESSE PERIODO
-- TEMOS UM CICLO DE 0.001s COM FREQUENCIA DE 1KHZ
--    __    __    __
-- __|  |__|  |__|  |
--
--|-----|     |--| 
-- 0.001s    0.0005s

-- O CLOCK DEVE INVERTER DUAS VEZES DENTRO DE UM PERIODO DE 0.001s
-- COMPONDO O NIVEL BAIXO POR 0.0005s E NIVEL ALTO PELO MESMO TEMPO


ENTITY CONVERSOR_1KHZ IS
PORT(
		CLK_I : IN STD_LOGIC;
		CLK_O : OUT STD_LOGIC
);
END CONVERSOR_1KHZ;

ARCHITECTURE LOGIC OF CONVERSOR_1KHZ IS
	SIGNAL SINAL_CLK : STD_LOGIC := '1';
BEGIN

PROCESS(CLK_I)
VARIABLE COUNT : INTEGER := 1;
BEGIN
	IF( CLK_I'EVENT AND CLK_I = '0') THEN

		COUNT := COUNT + 1;
		
		IF ( COUNT = 13500) THEN
		
			SINAL_CLK <= NOT SINAL_CLK;
			COUNT := 1;
			
		END IF;
	END IF;


END PROCESS;

CLK_O <= SINAL_CLK;


END LOGIC;