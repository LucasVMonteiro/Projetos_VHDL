library verilog;
use verilog.vl_types.all;
entity CONVERSOR_1KHZ_vlg_vec_tst is
end CONVERSOR_1KHZ_vlg_vec_tst;
