LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY BLOCO_PRINCIPAL IS 
PORT(
		CLOCK_IN : IN STD_LOGIC;
		SAIDA_R  : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
		SAIDA_G  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		
		);
END BLOCO_PRINCIPAL;

ARCHITECTURE LOGICA OF BLOCO_PRINCIPAL IS
--COMPONENTS



BEGIN



END LOGICA;
