LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-- ANODO COMUM
ENTITY DECODE_BCD_7SEG IS
	PORT(
			BCD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			OUT_7BIT : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
			);
END DECODE_BCD_7SEG;

ARCHITECTURE LOGICA OF DECODE_BCD_7SEG IS

BEGIN

WITH BCD SELECT  -- G F E D C B A --
	OUT_7BIT <= NOT "0111111" WHEN "0000",
					NOT "0000110" WHEN "0001",
					NOT "1011011" WHEN "0010",
					NOT "1001111" WHEN "0011",
					NOT "1100110" WHEN "0100",
					NOT "1101101" WHEN "0101",
					NOT "1111101" WHEN "0110",
					NOT "0000111" WHEN "0111",
					NOT "1111111" WHEN "1000",
					NOT "1101111" WHEN "1001",
					NOT "ZZZZZZZ" WHEN OTHERS;

END LOGICA;