library verilog;
use verilog.vl_types.all;
entity CONVERSOR_1KHZ_vlg_check_tst is
    port(
        CLK_O           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CONVERSOR_1KHZ_vlg_check_tst;
