LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BLOCO_PRINCIPAL IS 
PORT(
		CLOCK_IN : IN STD_LOGIC;
		
		TESTE_SINAL_FINAL_RED : OUT STD_LOGIC;
		TESTE_SINAL_FINAL_GREEN : OUT STD_LOGIC;
		TESTE_SINAL_CLKO_RED : OUT STD_LOGIC;
		TESTE_SINAL_CLKO_GREEN : OUT STD_LOGIC;
		TESTE_SINALTESTE_1SR : OUT STD_LOGIC;
		TESTE_SINALTESTE_1SG : OUT STD_LOGIC;
		
		SAIDA_R  : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
		SAIDA_G  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		
		
		);
END BLOCO_PRINCIPAL;

ARCHITECTURE LOGICA OF BLOCO_PRINCIPAL IS
--COMPONENTS

COMPONENT CONVERSOR_1KHZ IS
PORT(
		CLK_I : IN STD_LOGIC;
		CLK_O : OUT STD_LOGIC
);
END COMPONENT;

COMPONENT TEMPORIZADOR IS
PORT (
		CLK_I : IN STD_LOGIC;
		TEMPO : IN STD_LOGIC_VECTOR(4 DOWNTO 0); -- EM SEGUNDOS
		N_BITS : IN STD_LOGIC_VECTOR(4 DOWNTO 0); -- ATE 32 BITS
		CHIP_SELECT : IN STD_LOGIC;
		SINAL_FINAL : OUT STD_LOGIC;
		SINALTESTE_1S : OUT STD_LOGIC;
		CLK_O : OUT STD_LOGIC
);
END COMPONENT;

-- SIGNALS

SIGNAL SINAL_CLKO_CONVERSOR : STD_LOGIC;

SIGNAL SINAL_FINAL_RED : STD_LOGIC;
SIGNAL SINAL_CLKO_RED  : STD_LOGIC;

SIGNAL SINAL_FINAL_GREEN : STD_LOGIC;
SIGNAL SINAL_CLKO_GREEN  : STD_LOGIC;

SIGNAL BITS_RED : STD_LOGIC_VECTOR(17 DOWNTO 0):= "111111111111111111";
SIGNAL BITS_GREEN : STD_LOGIC_VECTOR(7 DOWNTO 0):= "00000000";

SIGNAL CHIP_SELECT : STD_LOGIC := '1';


BEGIN

CONVERSOR : CONVERSOR_1KHZ PORT MAP(CLOCK_IN,SINAL_CLKO_CONVERSOR);


TEMPORIZADOR_RED : TEMPORIZADOR PORT MAP(	
														SINAL_CLKO_CONVERSOR,
														"00101", -- 6  = 00110
														"10010", -- 18 = 10010
														'0',
														SINAL_FINAL_RED,
														TESTE_SINALTESTE_1SR,
														SINAL_CLKO_RED
														);
														
TEMPORIZADOR_GREEN : TEMPORIZADOR PORT MAP(	
															SINAL_CLKO_CONVERSOR,
															"00101", -- 6  = 00110
															"01000", -- 8  = 01000
															'1',
															SINAL_FINAL_GREEN,
															TESTE_SINALTESTE_1SG,
															SINAL_CLKO_GREEN
														);													
		TESTE_SINAL_FINAL_RED <= SINAL_FINAL_RED;
		TESTE_SINAL_FINAL_GREEN <= SINAL_FINAL_GREEN;
		TESTE_SINAL_CLKO_RED <= SINAL_CLKO_RED;
		TESTE_SINAL_CLKO_GREEN <= SINAL_CLKO_GREEN;
												
														
DESLOCADOR_RED:PROCESS(SINAL_CLKO_RED)

BEGIN
	IF(SINAL_CLKO_RED'EVENT AND SINAL_CLKO_RED = '0') THEN
		IF (BITS_RED = "000000000000000000") THEN
			BITS_RED <= "111111111111111111";
		END IF;
		IF (BITS_RED = "000000000000000001") THEN
			BITS_RED <= "000000000000000000";
		END IF;
		IF (BITS_RED > "000000000000000000") THEN
			BITS_RED <= STD_LOGIC_VECTOR( UNSIGNED(BITS_RED) / "000000000000000010");
		END IF;
	END IF;
END PROCESS DESLOCADOR_RED;

DESLOCADOR_GREEN:PROCESS(SINAL_CLKO_GREEN)

BEGIN
	IF(SINAL_CLKO_GREEN'EVENT AND SINAL_CLKO_GREEN = '0') THEN
		IF (BITS_GREEN = "00000000") THEN
			BITS_GREEN <= "11111111";
		END IF;
		IF (BITS_GREEN = "00000001") THEN
			BITS_GREEN <= "00000000";
		END IF;
		IF (BITS_GREEN > "00000000") THEN
			BITS_GREEN <= STD_LOGIC_VECTOR( UNSIGNED(BITS_GREEN) / "00000010");
		END IF;
	END IF;
END PROCESS DESLOCADOR_GREEN;

SAIDA_R <= BITS_RED;				
SAIDA_G <= BITS_GREEN;									
END LOGICA;
