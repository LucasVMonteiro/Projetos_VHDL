LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FSM_MEALY_2 IS
	PORT(
			X : IN STD_LOGIC;
			RST : IN STD_LOGIC;
			CLK : IN STD_LOGIC;
			y : OUT STD_LOGIC
			);
END FSM_MEALY_2;

ARCHITECTURE LOGIC OF FSM_MEALY_2 IS
	
-- SINAIS DO 1 FLIP FLOP D
	SIGNAL Q0 : STD_LOGIC := '0';
	SIGNAL D0 : STD_LOGIC := '0';
	
-- SINAIS DO 2 FLIP FLOP D
	SIGNAL Q1 : STD_LOGIC := '0';
	SIGNAL D1 : STD_LOGIC := '0';
	
	TYPE LIST_STATE IS( A, B, C);
	SIGNAL PR_STATE, NX_STATE: LIST_STATE;
	
BEGIN


	-- 	BLOCO COMBINACIONAL : PROCESSA
	-- O ESTADO ATUAL JUNTO A UMA ENTRADA
	-- E PRODUZ UMA SAIDA Y, E CALCULA O NX_STATE
	
	PROCESS( PR_STATE )
	BEGIN
	
		CASE PR_STATE IS
			WHEN A =>
				IF( X = '0' ) THEN
					Y <= '0';
					NX_STATE <= B;
				ELSE
					Y <= '0';
					NX_STATE <= A;
				END IF;
			
			WHEN B =>
				IF( X = '0' ) THEN
					Y <= '0';
					NX_STATE <= B;
				ELSE
					Y <= '0';
					NX_STATE <= C;
				END IF;		
			WHEN C =>
				IF( X = '0' ) THEN
					Y <= '1';
					NX_STATE <= A;
				ELSE
					Y <= '0';
					NX_STATE <= A;
				END IF;
			END CASE;
	END PROCESS;
	
		-- 	BLOCO SEQUENCIAL : CARREGA O PROXIMO
		-- ESTADO DENTRO DO ESTADO ATUAL
	
	PROCESS( CLK, RST )	
	BEGIN
		IF( RST = '1' ) THEN
			PR_STATE <= A;
		ELSIF( FALLING_EDGE(CLK)) THEN
			PR_STATE <= NX_STATE;
		END IF;
	END PROCESS;



END LOGIC;