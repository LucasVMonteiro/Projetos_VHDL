library verilog;
use verilog.vl_types.all;
entity BLOCO_CONTADOR23 is
    port(
        CLK_IN          : in     vl_logic;
        SAIDA           : out    vl_logic_vector(6 downto 0)
    );
end BLOCO_CONTADOR23;
