library verilog;
use verilog.vl_types.all;
entity BLOCO_CONTADOR59_vlg_check_tst is
    port(
        SAIDA           : in     vl_logic_vector(6 downto 0);
        sampler_rx      : in     vl_logic
    );
end BLOCO_CONTADOR59_vlg_check_tst;
