LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SEMAFORO IS 
PORT(
		CLK_IN : IN STD_LOGIC; -- CLOCK 50MHz
		SAIDA_R : OUT STD_LOGIC_VECTOR( 12 DOWNTO 0);
		SAIDA_G : OUT STD_LOGIC_VECTOR( 6 DOWNTO 0)
		
		);
END SEMAFORO;

ARCHITECTURE LOGIC OF SEMAFORO IS

SIGNAL LEDS_R : STD_LOGIC_VECTOR( 11 DOWNTO 0):= "111111111111";
SIGNAL LEDS_G : STD_LOGIC_VECTOR( 5 DOWNTO 0):= "000000";

SIGNAL LED_R  : STD_LOGIC := '1';
SIGNAL LED_G  : STD_LOGIC := '0';

CONSTANT TEMPO  : INTEGER := 6;
CONSTANT FREQUENCIA_CLK : INTEGER := 50000000;

BEGIN
SAIDA_R <= LED_R & LEDS_R;
SAIDA_G <= LED_G & LEDS_G;
PROCESS(CLK_IN)

	VARIABLE CONTADOR_CLK      : INTEGER := 1;
	--VARIABLE CONTADOR_SEGUNDOS : INTEGER := 1;
	VARIABLE TOGGLE : BIT := '0';

BEGIN

	IF( FALLING_EDGE(CLK_IN) ) THEN

		CONTADOR_CLK := CONTADOR_CLK + 1;
		
		IF( CONTADOR_CLK = FREQUENCIA_CLK ) THEN
			--CONTADOR_SEGUNDOS := CONTADOR_SEGUNDOS + 1;
			CONTADOR_CLK:=1;
			-- DESLOQUE 2 BITS RED A CADA 1 SEGUNDO
			IF(TOGGLE = '0') THEN
				
				IF( LEDS_R = "000000000000") THEN
					TOGGLE := '1';
					LEDS_G <= "111111";
					LED_R <= '0'; -- LED_R RECEBE 0
					LED_G <= '1';
				END IF;
				LEDS_R <= STD_LOGIC_VECTOR(SHIFT_RIGHT(UNSIGNED(LEDS_R),2));
		
			-- DESLOQUE 1 BIT A CADA 1 SEGUNDOS
			ELSIF( TOGGLE = '1') THEN
				
				IF( LEDS_G = "000000" ) THEN
					TOGGLE := '0';
					LEDS_R <= "111111111111";
					LED_R <= '1'; -- LED_R RECEBE 0
					LED_G <= '0';
				END IF;
				LEDS_G <= STD_LOGIC_VECTOR(SHIFT_RIGHT(UNSIGNED(LEDS_G),1));
			END IF;
			
			
		
		END IF;
		

	END IF;

END PROCESS;



END LOGIC;
