library verilog;
use verilog.vl_types.all;
entity BLOCO_CONTADOR59_vlg_vec_tst is
end BLOCO_CONTADOR59_vlg_vec_tst;
