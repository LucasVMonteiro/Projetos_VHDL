LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FSM_MEALY_1 IS
	PORT(
			X : IN STD_LOGIC;
			CLK : IN STD_LOGIC;
			y : OUT STD_LOGIC
			);
END FSM_MEALY_1;

ARCHITECTURE LOGIC OF FSM_MEALY_1 IS
	
-- SINAIS DO 1 FLIP FLOP D
	SIGNAL Q0 : STD_LOGIC := '0';
	SIGNAL D0 : STD_LOGIC := '0';
	
-- SINAIS DO 2 FLIP FLOP D
	SIGNAL Q1 : STD_LOGIC := '0';
	SIGNAL D1 : STD_LOGIC := '0';
	
	
	
BEGIN


	PROCESS( CLK )
		BEGIN
			IF( FALLING_EDGE(CLK) ) THEN
				Q0 <= D0;
				Q1 <= D1;
			END IF;
		END PROCESS;

	Y <= Q1 AND (NOT X);
	D1 <= Q0 AND X;
	D0 <= (NOT Q1) AND (NOT X);

END LOGIC;