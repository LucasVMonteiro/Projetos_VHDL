library verilog;
use verilog.vl_types.all;
entity BLOCO_CONTADOR23_vlg_vec_tst is
end BLOCO_CONTADOR23_vlg_vec_tst;
