library verilog;
use verilog.vl_types.all;
entity BLOCO_CONTADOR59_vlg_sample_tst is
    port(
        CLK_IN          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end BLOCO_CONTADOR59_vlg_sample_tst;
